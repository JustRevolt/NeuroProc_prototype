`define DATA_TYPE_SIZE 32

package types;
    typedef logic signed [`DATA_TYPE_SIZE-1:0] data_type;

endpackage
