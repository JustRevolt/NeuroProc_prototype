`define VIVADO_PRJ_USE
